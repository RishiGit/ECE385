module reg_8 (input  logic Clk, Reset, Load,
				  //Shift_In, Shift_En,
              input  logic [7:0]  D,
              //output logic Shift_Out,
              output logic [7:0]  Data_Out);

    always_ff @ (posedge Clk)
    begin
	 	 if (Reset) //notice, this is a sycnrhonous reset, which is recommended on the FPGA
			  Data_Out <= 8'h0;
		 else if (Load)
			  Data_Out <= D;
		 /*else if (Shift_En)
		 begin
			  //concatenate shifted in data to the previous left-most 3 bits
			  //note this works because we are in always_ff procedure block
			  Data_Out <= { Shift_In, Data_Out[7:1] }; 
	    end*/
    end
	
    //assign Shift_Out = Data_Out[0];

endmodule

module reg_4 (input  logic Clk, Reset, Load,
				  //Shift_In, Shift_En,
              input  logic [3:0]  D,
              //output logic Shift_Out,
              output logic [3:0]  Data_Out);

    always_ff @ (posedge Clk)
    begin
	 	 if (Reset) //notice, this is a sycnrhonous reset, which is recommended on the FPGA
			  Data_Out <= 4'h0;
		 else if (Load)
			  Data_Out <= D;
		 /*else if (Shift_En)
		 begin
			  //concatenate shifted in data to the previous left-most 3 bits
			  //note this works because we are in always_ff procedure block
			  Data_Out <= { Shift_In, Data_Out[3:1] }; 
	    end*/
    end
	
    //assign Shift_Out = Data_Out[0];

endmodule

module reg_16 (input logic Clk, Reset, Load,
				  //Shift_In, Shift_En,
              input  logic [15:0]  D,
              //output logic Shift_Out,
              output logic [15:0]  Data_Out);

    always_ff @ (posedge Clk)
    begin
	 	 if (Reset) //notice, this is a sycnrhonous reset, which is recommended on the FPGA
			  Data_Out <= 16'h0;
		 else if (Load)
			  Data_Out <= D;
		 /*else if (Shift_En)
		 begin
			  //concatenate shifted in data to the previous left-most 3 bits
			  //note this works because we are in always_ff procedure block
			  Data_Out <= { Shift_In, Data_Out[15:1] }; 
	    end*/
    end
	
    //assign Shift_Out = Data_Out[0];

endmodule

module reg_128 (input logic Clk, Reset, Load, first,
				  //Shift_In, Shift_En,
              input  logic [127:0]  D, d2,
              //output logic Shift_Out,
              output logic [127:0]  Data_Out);

    always_ff @ (posedge Clk)
    begin
		 if(first)
			Data_Out <= d2;
	 	 else if (Reset) //notice, this is a sycnrhonous reset, which is recommended on the FPGA
			  Data_Out <= 128'h0;
		 else if (Load)
			  Data_Out <= D;
		 /*else if (Shift_En)
		 begin
			  //concatenate shifted in data to the previous left-most 3 bits
			  //note this works because we are in always_ff procedure block
			  Data_Out <= { Shift_In, Data_Out[15:1] }; 
	    end*/
    end
	
    //assign Shift_Out = Data_Out[0];

endmodule

module eightreg_16 (input logic Clk, Reset, Load,
							input logic [15:0] D,
							input logic [2:0] SR1IN, SR2, DRIN,
							
							output logic [15:0] SR2O, SR1O);
		
		logic [7:0][15:0] regs;
		
		always_ff @ (posedge Clk)
		
			begin
					if(Reset)
						
						begin
						
							regs[0] <= 16'h0;
							regs[1] <= 16'h0;
							regs[2] <= 16'h0;
							regs[3] <= 16'h0;
							regs[4] <= 16'h0;
							regs[5] <= 16'h0;
							regs[6] <= 16'h0;
							regs[7] <= 16'h0;
							
					
						end
						
					else if (Load)
						
						case(DRIN)
							
								3'b000: regs[0] <= D;
								3'b001: regs[1] <= D;
								3'b010: regs[2] <= D;
								3'b011: regs[3] <= D;
								3'b100: regs[4] <= D;
								3'b101: regs[5] <= D;
								3'b110: regs[6] <= D;
								3'b111: regs[7] <= D;
								
								default ;
								
						endcase
						
			end
			
			always_comb
			
			begin
			
						case(SR1IN)
							
								3'b000: SR1O <= regs[0];
								3'b001: SR1O <= regs[1];
								3'b010: SR1O <= regs[2];
								3'b011: SR1O <= regs[3];
								3'b100: SR1O <= regs[4];
								3'b101: SR1O <= regs[5];
								3'b110: SR1O <= regs[6];
								3'b111: SR1O <= regs[7];
								
								default ;
								
						endcase
							
						case(SR2)
							
								3'b000: SR2O <= regs[0];
								3'b001: SR2O <= regs[1];
								3'b010: SR2O <= regs[2];
								3'b011: SR2O <= regs[3];
								3'b100: SR2O <= regs[4];
								3'b101: SR2O <= regs[5];
								3'b110: SR2O <= regs[6];
								3'b111: SR2O <= regs[7];
								
								default ;
								
						endcase
					
			end
		
endmodule	
							

module flip_flop (input  logic Clk, Reset, Load,
				  //Shift_In, Shift_En,
              input  logic  D,
              //output logic Shift_Out,
              output logic Data_Out);

    always_ff @ (posedge Clk)
    begin
	 	 if (Reset) //notice, this is a sycnrhonous reset, which is recommended on the FPGA
			  Data_Out <= 1'b0;
		 else if (Load)
			  Data_Out <= D;
		 /*else if (Shift_En)
		 begin
			  //concatenate shifted in data to the previous left-most 3 bits
			  //note this works because we are in always_ff procedure block
			  Data_Out <= { Shift_In, Data_Out[15:1] }; 
	    end*/
    end
	
    //assign Shift_Out = Data_Out[0];

endmodule
